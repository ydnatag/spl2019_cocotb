--------------------------------------------------------------------------------
-- Company: Satellogic S.A
--
-- File: axi_lite_slave_int.vhdl
-- Description: 
--
-- AXI Lite Slave Interface for any ip core. Based in Xilinx automagic core.
--
-- Author: Xilinx, David Caruso
--
--------------------------------------------------------------------------------

entity example is
    generic ();
    port ();
end example;

architecture rtl of example is
end rtl;
