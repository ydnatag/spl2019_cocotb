
module example();
endmodule
