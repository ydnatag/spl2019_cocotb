`timescale 1ns/1ps
module example();
endmodule
